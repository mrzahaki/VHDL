-- W T A
--library IEEE;
--use IEEE.STD_LOGIC_1164.all;

package std_type is

--TYPE integer_vector	is array(NATURAL range<>) of INTEGER;
  TYPE boolean_vector	is array(NATURAL range<>) of BOOLEAN;--vhdl 2008
  TYPE integer_vector	is array(NATURAL range<>) of INTEGER;


end package std_type;
PACKAGE BODY std_type IS
END PACKAGE BODY std_type;
